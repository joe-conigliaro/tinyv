// Copyright (c) 2020-2023 Joe Conigliaro. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module ast

import tinyv.token

// NOTE: this is just a very naive example of how it could possibly work.
// actual implementation may work during AST -> IR (or not). it may also
// need type information which we don't have here. as I said, just an example.
pub fn(m &MatchExpr) desugar() Expr {
	mut if_expr := ast.IfExpr{}
	for i, branch in m.branches {
		mut branch_cond := empty_expr
		for cond in branch.cond {
			op := if cond in [ast.Ident, ast.SelectorExpr] { token.Token.key_is } else { token.Token.eq }
			c := ast.InfixExpr{lhs: m.expr, op: op, rhs: cond}
			if branch_cond !is EmptyExpr {
				branch_cond = InfixExpr{lhs: branch_cond, op: .logical_or, rhs: c}
			} else {
				branch_cond = c
			}
		}
		if_expr2 := ast.IfExpr{
			cond: branch_cond
			stmts: branch.stmts
		}
		if i == 0 {
			if_expr = if_expr2
		} else {
			if_expr = ast.IfExpr{...if_expr else_expr: if_expr2}
		}
	}
	return if_expr
}