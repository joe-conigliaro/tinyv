module main

fn main() {
    a, b := 1, 2
	arr1 := [1,2,3,4]
	// arr2 := []string{len: 2, cap :2} // TODO: see comment in parser
	arr2 := []string{len: 2}
	x := foo[1]()

}
