module types

pub type Object = Number | Struct

pub struct Type{
	object Object
}

struct Number{

}

struct Struct{

}