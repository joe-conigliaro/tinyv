module types

const(
	// universe = &Scope
)