module pref

pub struct Preferences {
pub:
	verbose bool
}
