module types

struct Checker {

}

pub fn new_checker() &Checker {
	return &Checker{

	}
}
