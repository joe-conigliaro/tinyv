module main

fn main() {
    a, b := 1, 2

    x := foo[1]()
}