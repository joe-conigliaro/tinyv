module pref

pub struct Preferences {
pub:
	debug   bool
	verbose bool
}
